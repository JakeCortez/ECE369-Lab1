`timescale 1ns / 1ps

module InstructionFetchUnit_tb()


endmodule